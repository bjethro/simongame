`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 02/25/2016 12:41:21 PM
// Design Name:
// Module Name: Checking_nbits
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
// Check if one-bit input is correct
module Checking_1bit(
    output          correct,
    output [1:0]    led_pressed,
    input           clock,
    input           right_pressed,
    input           left_pressed,
    input           enable,
    input           bit_gen      // bit generated by random number generator
    );

reg         correct_reg;
reg  [1:0]  led_pressed_reg;

assign      correct         = correct_reg;
assign      led_pressed     = led_pressed_reg;

always @(posedge clock) begin
    if (enable) begin
        if (right_pressed == 1) begin
            led_pressed_reg     <= 0'b01;
            if (bit_gen == 1)   correct_reg <= 1;
            else                correct_reg <= 0;
            end
        else if (left_pressed == 1) begin
            led_pressed_reg     <= 0'b10;
            if (bit_gen == 0)   correct_reg <= 1;
            else                correct_reg <= 0;
            end
        else    led_pressed_reg <= 0'b00;
        end
    else
        led_pressed_reg         <= 0'b00;
    end

endmodule
